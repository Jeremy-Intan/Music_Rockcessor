module wb_stage();

input wire [15:0] rd_data;
input wire [3:0] rd_addr;
input wire [15:0] bd_data;
input wire [16:0] n_mem_data;
input wire [1535:0] b_mem_data;


endmodule
