module dec_stage();



endmodule
