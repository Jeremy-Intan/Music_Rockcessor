module cmpalu(input clk, input start, input [63:0] bitcolumn, input [23:0] bitrowtop, input [23:0] bitrowbot, input nextrowtopready, input nextrowbotready, input nextcolumnready, input lastcolumn, output [15:0] result, output done, output nextcolumn, output nextrowtop, output nextrowbot);

//Takes in slices of a 64x24 bitmap and determines how far it should be shifted left and down, and whether or not it should be scaled by 2x

//output signals
reg finished;
reg botrowchecked;
reg toprowchecked;
assign done = finished;
assign nextrowtop = toprowchecked;
assign nextrowbot = botrowchecked;

//[4:0] = lshift
//[10:5] = dshift
//[11] = scale 2x horizontal
//[12] = scale 2x vertical
reg [15:0] res;
assign result = res;

//input
//bitmap staging
reg [63:0] currcol;
reg [23:0] currrowtop;
reg [23:0] currrowbot;

//number of empty columns and rows
reg [4:0] emptycolumns;
reg [5:0] emptyrows;
reg [5:0] emptyrowsupper;
reg [5:0] emptyrowslower;

//booleans

//1 indicates that the row or column needs to be checked
reg checkcol;
reg checkrowtop;
reg checkrowbot;

//1 indicates that the boundary has been found
reg lboundaryfound;
reg topboundaryfound;
reg botboundaryfound;

//1 indicates that the boundary has been stored in the result
reg lboundarystored;
reg topboundarystored;
reg botboundarystored;

//[0] is the calculation for left columns
//[1] is the calculation for bot rows
//[2] is the calculation for horizontal scaling
//[3] is the calculation for vertical scaling
reg [3:0] calcdone;

//Row check logic
//checks from top to bot
//and bot to top

//finds empty rows on top
always @(posedge clk) begin
    casez ({checkrowtop, currrowtop})
        //check each row only once
        //checkrow, rowempty
        {1'b1,24'h00} : begin
                        emptyrowsupper <= emptyrowsupper + 1;
                        checkrowtop <= 1'b0;
                        toprowchecked <= 1'b1;
                        end

        //don't cares if we shouldn't check row
        {1'b1, 24'h??} : emptyrowsupper <= emptyrowsupper;

        //checkrow, row not empty
        default :   begin
                    emptyrowsupper <= emptyrowsupper;
                    topboundaryfound <= 1'b1;
                    checkrowtop <= 1'b0;
                    toprowchecked <= 1'b1;
                    end
    endcase
end

//finds empty rows on bot
always @(posedge clk) begin
    casez ({checkrowbot, currrowbot})
        //check each row only once
        //checkrow, rowempty
        {1'b1,24'h00} : begin
                        emptyrowslower <= emptyrowslower + 1;
                        checkrowbot <= 1'b0;
                        botrowchecked <= 1'b1;
                        end

        //don't cares if we shouldn't check row
        {1'b1, 24'h??} : emptyrowslower <= emptyrowslower;

        //checkrow, row not empty
        default :   begin
                    emptyrowslower <= emptyrowslower;
                    botboundaryfound <= 1'b1;
                    checkrowbot <= 1'b0;
                    botrowchecked <= 1'b1;
                    end
    endcase
end

//row store logic
always @(posedge clk) begin
    
    //store number of empty rows top
    case ({topboundaryfound, topboundarystored})
        2'b10 : begin
                emptyrows <= emptyrows + emptyrowsupper;
                topboundarystored <= 1'b1;
                end
        default: emptyrows <= emptyrows;
    endcase

    //store number of empty rows bot
    case ({botboundaryfound, botboundarystored})
        2'b10 : begin
                emptyrows <= emptyrows + emptyrowslower;
                res [10:5] <= emptyrowslower;
                calcdone[2] <= 1'b1;
                botboundarystored <= 1'b1;
                end 
        default : emptyrows <= emptyrows;
    endcase

    case ({topboundarystored, botboundarystored, emptyrows[5]})
        //row calcs done, check if num empty rows >= 32
        3'b111 :    begin
                    res [12] <= 1'b1;
                    calcdone[3] <= 1'b1;
                    end
        3'b110 :    begin
                    res [12] <= 1'b0;
                    calcdone[3] <= 1'b1;
                    end
        default:    res[12] <= res[12];
    endcase
end

//Column check logic
always @(posedge clk) begin
    case ({lboundaryfound, lboundarystored})
    //store lshift in result once first boundary has been found
        2'b10 :  begin
                res [5:0] <= emptycolumns;
                calcdone [0] <= 1'b1;
                end
        default : emptycolumns <= emptycolumns;
    endcase

    case ({lastcolumn, emptycolumns[4]})
        //last column, 12 or greater empty columns
        //presently checks for 16 or greater, update later
        2'b11 :    begin 
                    res [11] <= 1'b1;
                    calcdone [1] <= 1'b1;
                    end
        2'b10 :     begin
                    res [11] <= 1'b0;
                    calcdone [1] <= 1'b1;
                    end
        default : calcdone[1] <= calcdone[1];
    endcase
end

always @(posedge clk) begin

    casez ({checkcol, currcol})
        //check each column only once
        //checkcolumn, column empty
        65'h10000 : begin
                    emptycolumns <= emptycolumns + 1;
                    checkcol <= 1'b0;
                    end

        //don't cares if column has been checked
        65'h0????:  begin
                    emptycolumns <= emptycolumns;
                    end

        //checkcolumn, column not empty
        default :   begin
                    emptycolumns <= emptycolumns;
                    checkcol <= 1'b0;
                    lboundaryfound <= 1'b1;
                    end
    endcase
end

//move current row and column into reg banks
always @(posedge clk)  begin
    //next column
    case (nextcolumnready)
        1'b1  : begin
                currcol <= bitcolumn;
                checkcol <= 1'b1;
                end
        default: currcol <= currcol;
    endcase  

    //nexttoprow
    case (nextrowtopready)
        1'b1  : begin
                currrowtop <= bitrowtop;
                checkrowtop <= 1'b1;
                end
        default: currrowtop <= currrowtop;
    endcase

    //nextbotrow
    case (nextrowbotready)
        1'b1  : begin
                currrowbot <= bitrowbot;
                checkrowbot <= 1'b1;
                end
        default: currrowbot <= currrowbot;
    endcase  

    //once all 4 calcs are done, send finish signal
    case (calcdone)
        4'b1111 : finished <= 1'b1; 
        default : finished <= 1'b0;
    endcase

    //reset alu on start
    case (start)
        1'b1 : begin
                emptycolumns <= 5'b0;
                emptyrows <= 6'b0;
                emptyrowsupper <= 6'b0;
                emptyrowslower <= 6'b0;
                lboundaryfound <= 1'b0;
                lboundarystored <= 1'b0;
                topboundaryfound <= 1'b0;
                botboundaryfound <= 1'b0;
                topboundarystored <= 1'b0;
                botboundarystored <= 1'b0;
                res <= 16'h0;
				calcdone<= 4'b0;
                end
        default : finished <= 1'b0;
    endcase
end

endmodule
        