module inst_stage();



endmodule
