module wb_stage();



endmodule
