
module audio_clk (
	audio_clk_clk,
	ref_clk_clk,
	ref_reset_reset,
	reset_source_reset);	

	output		audio_clk_clk;
	input		ref_clk_clk;
	input		ref_reset_reset;
	output		reset_source_reset;
endmodule
