module inst_tb();

reg clk, rst_n;
reg stall;
reg [15:0] branch_pc;
reg branch_to_new;
wire [15:0] pc;
wire [15:0] inst;
wire inst_invalid;

inst_stage iDUT(.clk(clk), .rst_n(rst_n), .stall(stall), .branch_pc(branch_pc), .branch_to_new(branch_to_new), .pc(pc), .inst(inst), .inst_invalid(inst_invalid));

initial begin
clk = 0;
rst_n = 0;
stall = 0;
branch_pc = 0;
branch_to_new = 0;
@(negedge clk);
rst_n = 1;
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
branch_pc = 3;
branch_to_new = 1;
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
branch_to_new = 0;
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
branch_pc = 3;
branch_to_new = 0;
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
branch_pc = 9;
branch_to_new = 1;
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
branch_to_new = 0;
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
branch_pc = 12;
branch_to_new = 1;
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
branch_to_new = 0;
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
stall = 1;
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
@(posedge clk);
@(negedge clk);
$display("pc %d, inst %b, inst_invalid %b", pc, inst, inst_invalid);
$stop;
end


always begin
#2 clk = ~clk;
end

endmodule
